library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- X,Y to Relative X,Y
entity ExplosionLogic is
	Port ( 	Clk : in STD_LOGIC;
			X : in INTEGER;
			Y : in INTEGER;
			staticWallPresent : in STD_LOGIC;
			breakableWallPresent : in STD_LOGIC;
			bombExploding : in STD_LOGIC;
			explosionPresent : out STD_LOGIC ); -- Whether an explosion is present here
end ExplosionLogic;

architecture Behavioral of ExplosionLogic is
type matrix is array(0 to 28, 0 to 38) of STD_LOGIC_VECTOR ( 0 to 5 );
signal explosionLocation : matrix := (
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000"),
									("000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000","000000")
								);
begin
	process(Clk)
	variable matrixX : INTEGER;
	variable matrixY : INTEGER;
	variable neightbourExpl : STD_LOGIC; -- Tell if for the current iteration, there is a neightboor with an explosion
	begin
		If( Clk'Event and Clk = '1' ) then
			-- Compute the matrixX and matrixY
			If ((X >= 8 and Y >= 8 ) and (X < (640-8) and Y < (480-8) )) then
				matrixX := (((Y+8)/16)-1);
				matrixY := (((X+8)/16)-1);
				-- First, check if there is a bomb and plant it
				If (bombExploding = '1') then
					explosionLocation(matrixX, matrixY) <= "111111"; -- This is a bomb
				End If;
				-- Second, remove a already implemented bomb if it's not present anymore
				If (explosionLocation(matrixX, matrixY) = "111111") and bombExploding = '0' then
					explosionLocation(matrixX, matrixY) <= "000000";
				End If;
				-- Third, update current grid according to neightboors, (only update distance if not already explosion)
				neightbourExpl := '0'; -- If we go into no If, there is no neightboor with an explosion
				-- Explosion from up
				If (matrixX > 0) then
					If (explosionLocation(matrixX - 1, matrixY)(0) = '1' and explosionLocation(matrixX - 1, matrixY)(4 to 5) /= "00") then -- There is an explosion from top
						neightbourExpl := '1';
						explosionLocation(matrixX, matrixY) (0 to 3) <= "1000";
						If (explosionLocation(matrixX, matrixY) (4 to 5) = "00") then -- This is the first time we update the distance
							If (explosionLocation(matrixX - 1, matrixY)(4 to 5) = "11") then
								explosionLocation(matrixX, matrixY) (4 to 5) <= "10";
							End If;
							If (explosionLocation(matrixX - 1, matrixY)(4 to 5) = "10") then
								explosionLocation(matrixX, matrixY) (4 to 5) <= "01";
							End If;
							If (explosionLocation(matrixX - 1, matrixY)(4 to 5) = "01") then
								explosionLocation(matrixX, matrixY) (4 to 5) <= "00";
							End If;
						End If;
					End If;
				End If;
				-- Explosion from right
				If (matrixY < 38) then
					If (explosionLocation(matrixX, matrixY + 1)(1) = '1' and explosionLocation(matrixX, matrixY + 1)(4 to 5) /= "00") then -- There is an explosion from right
						neightbourExpl := '1';
						explosionLocation(matrixX, matrixY) (0 to 3) <= "0100";
						If (explosionLocation(matrixX, matrixY) (4 to 5) = "00") then -- This is the first time we update the distance
							If (explosionLocation(matrixX, matrixY + 1)(4 to 5) = "11") then
								explosionLocation(matrixX, matrixY) (4 to 5) <= "10";
							End If;
							If (explosionLocation(matrixX, matrixY + 1)(4 to 5) = "10") then
								explosionLocation(matrixX, matrixY) (4 to 5) <= "01";
							End If;
							If (explosionLocation(matrixX, matrixY + 1)(4 to 5) = "01") then
								explosionLocation(matrixX, matrixY) (4 to 5) <= "00";
							End If;
						End If;
					End If;
				End If;
				-- Explosion from down
				If (matrixX < 28) then
					If (explosionLocation(matrixX + 1, matrixY)(2) = '1' and explosionLocation(matrixX + 1, matrixY)(4 to 5) /= "00") then -- There is an explosion from down
						neightbourExpl := '1';
						explosionLocation(matrixX, matrixY) (0 to 3) <= "0010";
						If (explosionLocation(matrixX, matrixY) (4 to 5) = "00") then -- This is the first time we update the distance
							If (explosionLocation(matrixX + 1, matrixY)(4 to 5) = "11") then
								explosionLocation(matrixX, matrixY) (4 to 5) <= "10";
							End If;
							If (explosionLocation(matrixX + 1, matrixY)(4 to 5) = "10") then
								explosionLocation(matrixX, matrixY) (4 to 5) <= "01";
							End If;
							If (explosionLocation(matrixX + 1, matrixY)(4 to 5) = "01") then
								explosionLocation(matrixX, matrixY) (4 to 5) <= "00";
							End If;
						End If;
					End If;
				End If;
				-- Explosion from left
				If (matrixY > 0) then
					If (explosionLocation(matrixX, matrixY - 1)(3) = '1' and explosionLocation(matrixX, matrixY - 1)(4 to 5) /= "00") then -- There is an explosion from left
						neightbourExpl := '1';
						explosionLocation(matrixX, matrixY) (0 to 3) <= "0001";
						If (explosionLocation(matrixX, matrixY) (4 to 5) = "00") then -- This is the first time we update the distance
							If (explosionLocation(matrixX, matrixY - 1)(4 to 5) <= "11") then
								explosionLocation(matrixX, matrixY) (4 to 5) <= "10";
							End If;
							If (explosionLocation(matrixX, matrixY - 1)(4 to 5) = "10") then
								explosionLocation(matrixX, matrixY) (4 to 5) <= "01";
							End If;
							If (explosionLocation(matrixX, matrixY - 1)(4 to 5) = "01") then
								explosionLocation(matrixX, matrixY) (4 to 5) <= "00";
							End If;
						End If;
					End If;
				End If;
				-- If there was no neighbour detected, remove the explosion
				If (neightbourExpl = '0') then
					explosionLocation(matrixX, matrixY) <= "000000";
				End If;
				-- Fourth, tell whether there is an explosion
				If (explosionLocation(matrixX, matrixY) /= "000000") then
					explosionPresent <= '1';
				Else
					explosionPresent <= '0';
				End If;
			End If;
		End if;
	end process; 
end Behavioral;