library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Animated Sprite
-- animationSeq:
-- 1 : Down Idle
-- 2 : Down Move1
-- 3 : Down Move2
-- 11 : Left Idle
-- 12 : Left Move1
-- 13 : Left Move2
-- 21 : Up Idle
-- 22 : Up Move1
-- 23 : Up Move2
-- 31 : Right Idle
-- 32 : Right Move1
-- 33 : Right Move2

entity CharacterAnimatedSprite is
    Port ( relativeX : in INTEGER;
           relativeY : in INTEGER;
		   drawIt : in STD_LOGIC;
		   animationSeq : in INTEGER;
		   RGB : out STD_LOGIC_VECTOR (0 to 2) );
end CharacterAnimatedSprite;

architecture Behavioral of CharacterAnimatedSprite is
begin
	-- Begin of Animated Sprite Code
	-- From char_down_idle.png
	RGB <= 	"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 3) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 4) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 4) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 4) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 5) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 5) and (relativeY = 5)) else
			"100" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 5) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 5) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 5) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 5) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 5) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 5) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 6) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 6) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 6) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 6) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 6) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 6) and (relativeY = 13)) else
			"100" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 7) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 7) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 7) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 7) and (relativeY = 5)) else
			"100" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 7) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 7) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 7) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 7) and (relativeY = 9)) else
			"110" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 7) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 7) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 8) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 8) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 8) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 8) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 8) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 8) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 9) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 9) and (relativeY = 5)) else
			"100" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 9) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 9) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 9) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 9) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 9) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 9) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 10) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 10) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 10) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 1) and (relativeX = 11) and (relativeY = 11)) else
	-- End of Sprite Code
	-- From char_down_move1.png
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 4) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 4) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 5) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 5) and (relativeY = 5)) else
			"100" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 5) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 5) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 5) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 5) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 5) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 6) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 6) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 6) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 6) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 6) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 7) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 7) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 7) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 7) and (relativeY = 5)) else
			"100" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 7) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 7) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 7) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 7) and (relativeY = 9)) else
			"110" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 7) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 8) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 8) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 8) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 8) and (relativeY = 9)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 8) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 8) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 9) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 9) and (relativeY = 5)) else
			"100" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 9) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 9) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 9) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 9) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 9) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 9) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 9) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 10) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 10) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 2) and (relativeX = 10) and (relativeY = 13)) else
	-- End of Sprite Code
	-- From char_down_move2.png
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 4) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 4) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 4) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 5) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 5) and (relativeY = 5)) else
			"100" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 5) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 5) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 5) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 5) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 5) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 5) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 5) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 6) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 6) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 6) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 6) and (relativeY = 9)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 6) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 6) and (relativeY = 13)) else
			"100" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 7) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 7) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 7) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 7) and (relativeY = 5)) else
			"100" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 7) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 7) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 7) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 7) and (relativeY = 9)) else
			"110" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 7) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 8) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 8) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 8) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 8) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 8) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 9) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 9) and (relativeY = 5)) else
			"100" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 9) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 9) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 9) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 9) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 9) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 10) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 3) and (relativeX = 10) and (relativeY = 11)) else
	-- End of Sprite Code
	-- From char_left_idle.png
			"100" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 4) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 5) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 5) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 5) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 5) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 5) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 5) and (relativeY = 7)) else
			"001" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 5) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 6) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 6) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 6) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 6) and (relativeY = 9)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 6) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 6) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 7) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 7) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 7) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 7) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 7) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 7) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 7) and (relativeY = 9)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 7) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 7) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 7) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 8) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 8) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 8) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 8) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 8) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 8) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 8) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 8) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 8) and (relativeY = 13)) else
			"100" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 9) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 9) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 9) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 9) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 9) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 9) and (relativeY = 7)) else
			"001" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 9) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 9) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 10) and (relativeY = 2)) else
			"100" when ((drawIt = '1') and (animationSeq = 11) and (relativeX = 10) and (relativeY = 3)) else
	-- End of Sprite Code
	-- From char_left_move1.png
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 5) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 5) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 5) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 5) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 5) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 5) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 5) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 5) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 6) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 6) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 6) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 6) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 6) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 6) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 7) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 7) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 7) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 7) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 7) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 7) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 7) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 7) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 8) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 8) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 8) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 8) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 8) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 8) and (relativeY = 8)) else
			"001" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 8) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 8) and (relativeY = 13)) else
			"100" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 9) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 9) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 9) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 9) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 9) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 9) and (relativeY = 8)) else
			"001" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 9) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 9) and (relativeY = 13)) else
			"100" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 10) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 10) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 10) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 12) and (relativeX = 10) and (relativeY = 13)) else
	-- End of Sprite Code
	-- From char_left_move2.png
			"100" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 4) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 5) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 5) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 5) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 5) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 5) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 5) and (relativeY = 8)) else
			"001" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 5) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 5) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 5) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 6) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 6) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 6) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 6) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 6) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 7) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 7) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 7) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 7) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 7) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 7) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 7) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 8) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 8) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 8) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 8) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 8) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 8) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 8) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 8) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 8) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 9) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 9) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 9) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 9) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 9) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 9) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 9) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 9) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 10) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 13) and (relativeX = 10) and (relativeY = 4)) else
	-- End of Sprite Code
	-- From char_up_idle.png
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 3) and (relativeY = 8)) else
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 3) and (relativeY = 9)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 4) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 5) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 5) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 5) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 5) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 5) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 5) and (relativeY = 7)) else
			"001" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 5) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 5) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 6) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 6) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 6) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 6) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 6) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 6) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 6) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 6) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 6) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 7) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 7) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 7) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 7) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 7) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 7) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 7) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 7) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 8) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 8) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 8) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 8) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 8) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 8) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 8) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 8) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 8) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 9) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 9) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 9) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 9) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 9) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 9) and (relativeY = 7)) else
			"001" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 9) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 9) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 10) and (relativeY = 8)) else
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 11) and (relativeY = 8)) else
			"100" when ((drawIt = '1') and (animationSeq = 21) and (relativeX = 11) and (relativeY = 9)) else
	-- End of Sprite Code
	-- From char_up_move1.png
			"100" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 3) and (relativeY = 9)) else
			"100" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 3) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 4) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 4) and (relativeY = 9)) else
			"100" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 4) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 5) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 5) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 5) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 5) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 5) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 5) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 6) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 6) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 6) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 6) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 6) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 6) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 6) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 6) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 7) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 7) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 7) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 7) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 7) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 7) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 7) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 7) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 8) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 8) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 8) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 8) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 8) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 8) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 8) and (relativeY = 9)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 8) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 8) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 9) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 9) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 9) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 9) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 9) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 9) and (relativeY = 7)) else
			"001" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 9) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 9) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 9) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 10) and (relativeY = 8)) else
			"100" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 10) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 22) and (relativeX = 10) and (relativeY = 12)) else
	-- End of Sprite Code
	-- From char_up_move2.png
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 4) and (relativeY = 8)) else
			"100" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 4) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 4) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 5) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 5) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 5) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 5) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 5) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 5) and (relativeY = 7)) else
			"001" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 5) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 5) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 5) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 6) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 6) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 6) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 6) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 6) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 6) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 6) and (relativeY = 9)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 6) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 6) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 7) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 7) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 7) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 7) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 7) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 7) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 7) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 7) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 8) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 8) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 8) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 8) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 8) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 8) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 8) and (relativeY = 9)) else
			"001" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 8) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 9) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 9) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 9) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 9) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 9) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 9) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 10) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 10) and (relativeY = 9)) else
			"100" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 10) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 11) and (relativeY = 9)) else
			"100" when ((drawIt = '1') and (animationSeq = 23) and (relativeX = 11) and (relativeY = 10)) else
	-- End of Sprite Code
	-- From char_right_idle.png
			"100" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 5) and (relativeY = 2)) else
			"100" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 5) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 6) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 6) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 6) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 6) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 6) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 6) and (relativeY = 7)) else
			"001" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 6) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 6) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 7) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 7) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 7) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 7) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 7) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 7) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 7) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 7) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 7) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 8) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 8) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 8) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 8) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 8) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 8) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 8) and (relativeY = 9)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 8) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 8) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 8) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 9) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 9) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 9) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 9) and (relativeY = 9)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 9) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 9) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 10) and (relativeY = 2)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 10) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 10) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 10) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 10) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 10) and (relativeY = 7)) else
			"001" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 10) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 31) and (relativeX = 11) and (relativeY = 12)) else
	-- End of Sprite Code
	-- From char_right_move1.png
			"100" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 5) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 5) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 5) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 5) and (relativeY = 13)) else
			"100" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 6) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 6) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 6) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 6) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 6) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 6) and (relativeY = 8)) else
			"001" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 6) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 6) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 7) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 7) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 7) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 7) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 7) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 7) and (relativeY = 8)) else
			"001" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 7) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 7) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 8) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 8) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 8) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 8) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 8) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 8) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 8) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 8) and (relativeY = 11)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 9) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 9) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 9) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 9) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 9) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 9) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 10) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 10) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 10) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 10) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 10) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 10) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 10) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 32) and (relativeX = 10) and (relativeY = 12)) else
	-- End of Sprite Code
	-- From char_right_move2.png
			"100" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 5) and (relativeY = 3)) else
			"100" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 5) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 6) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 6) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 6) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 6) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 6) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 6) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 6) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 6) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 7) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 7) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 7) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 7) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 7) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 7) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 7) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 7) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 7) and (relativeY = 12)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 8) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 8) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 8) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 8) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 8) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 8) and (relativeY = 8)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 8) and (relativeY = 10)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 9) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 9) and (relativeY = 4)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 9) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 9) and (relativeY = 10)) else
			"100" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 9) and (relativeY = 13)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 10) and (relativeY = 3)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 10) and (relativeY = 4)) else
			"100" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 10) and (relativeY = 5)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 10) and (relativeY = 6)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 10) and (relativeY = 7)) else
			"111" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 10) and (relativeY = 8)) else
			"001" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 10) and (relativeY = 11)) else
			"100" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 10) and (relativeY = 12)) else
			"100" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 10) and (relativeY = 13)) else
			"100" when ((drawIt = '1') and (animationSeq = 33) and (relativeX = 11) and (relativeY = 12)) else
			"000";
	-- End of Sprite Code
end Behavioral;