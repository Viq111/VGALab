library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- X,Y to Relative X,Y
entity DestructibleWallLocalCoordinates is
	Port ( 	Clk : in STD_LOGIC;
			X : in INTEGER;
			Y : in INTEGER;
			relativeX : out INTEGER;
			relativeY : out INTEGER;
			drawIt : out STD_LOGIC );
end DestructibleWallLocalCoordinates;

architecture Behavioral of DestructibleWallLocalCoordinates is

type matrix is array(0 to 28, 0 to 38) of STD_LOGIC;
signal WallLocation : matrix := (	
									"010100000000000000000000000000000000001",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"000000000000000000000000000000000000000",
									"100000000000000000000000000000000000001"
								);

begin
	--drawIt <= '1' when ((WallLocation((((X+8)/16)-1), (((Y+8)/16)-1)) = '1') and ((X >= 8 and Y >= 8 ) or (X <= (640-8) and Y <= (480-8) ))) else '0';
	relativeX <= (X+8) mod 16;
	relativeY <= (Y+8) mod 16;
	process(Clk)
	begin
		if( Clk'Event and Clk = '1' ) then
			If ((X >= 8 and Y >= 8 ) and (X <= (640-8) and Y <= (480-8) )) then
				If WallLocation((((Y+8)/16)-1), (((X+8)/16)-1)) = '1' then
					drawIt <= '1';
				Else
					drawIt <= '0';
				End If;
			Else
				drawIt <= '0';
			End If;
		end if;
	end process; 
end Behavioral;