library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- X,Y to Relative X,Y
entity DestructibleWallLocalCoordinates is
	Port ( 	Clk : in STD_LOGIC;
			X : in INTEGER;
			Y : in INTEGER;
			relativeX : out INTEGER;
			relativeY : out INTEGER;
			drawIt : out STD_LOGIC;
			Interact : in STD_LOGIC	);
end DestructibleWallLocalCoordinates;

architecture Behavioral of DestructibleWallLocalCoordinates is

type matrix is array(0 to 28, 0 to 38) of STD_LOGIC;
signal WallLocation : matrix := (	
								"000000101000010010000010000000000100000",
								"001010000000000000000000000000000000001",
								"100010010000000000000010000010000000000",
								"000000000000000000000000000000100000100",
								"010000100100010010000100001000001000000",
								"000000000000000000000000000000000000001",
								"010010000000000000010100000101000000001",
								"000000001000100010000000000000000000000",
								"001000100000000000100000010001000100000",
								"000000001000001000000000100000000000001",
								"000000000001000000010000000000000000000",
								"000000000000000000000000001000000000000",
								"100100000000100001000001000000100001000",
								"000000000000000000001000000000000000001",
								"001001000100000001000000000100001001000",
								"000000000000000000000000100000000000000",
								"101000000000100000000000000001000000010",
								"000010000000000000000000000000001000000",
								"000000000010000010000000100100000000101",
								"001000000000000000100000000000000000000",
								"000000001000000100001000000000100001001",
								"000000000000000000100000101000000000000",
								"001001000010001000000100000001010010000",
								"000010000000000000000000001000000000101",
								"100000000010010000000101000000010010000",
								"001000000000000000100000000000000000001",
								"100000000001000010001000000000000000100",
								"000010000000001000100010000000000000000",
								"101000000001000000000000000000001001000"
								);

begin
	--drawIt <= '1' when ((WallLocation((((X+8)/16)-1), (((Y+8)/16)-1)) = '1') and ((X >= 8 and Y >= 8 ) or (X <= (640-8) and Y <= (480-8) ))) else '0';
	relativeX <= (X+8) mod 16;
	relativeY <= (Y+8) mod 16;
	process(Clk)
	begin
		if( Clk'Event and Clk = '1' ) then
			-- Draw Breakable Wall
			If ((X >= 8 and Y >= 8 ) and (X < (640-8) and Y < (480-8) )) then
				If WallLocation((((Y+8)/16)-1), (((X+8)/16)-1)) = '1' then
					drawIt <= '1';
				Else
					drawIt <= '0';
				End If;
			Else
				drawIt <= '0';
			End If;
			
			-- Destroy
			If ((X >= 8 and Y >= 8 ) and (X < (640-8) and Y < (480-8) )) then
				If (WallLocation((((Y+8)/16)-1), (((X+8)/16)-1)) = '1' and Interact = '1') then
					WallLocation((((Y+8)/16)-1), (((X+8)/16)-1)) <= '0';
				End If;
			End If;
		end if;
	end process; 
end Behavioral;